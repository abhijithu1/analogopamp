magic
tech sky130A
magscale 1 2
timestamp 1742637551
<< error_s >>
rect -978 -336 -920 -330
rect -978 -370 -966 -336
rect -978 -376 -920 -370
rect -978 -548 -920 -542
rect -978 -582 -966 -548
rect -978 -588 -920 -582
rect -1518 -1116 -1460 -1110
rect -518 -1116 -460 -1110
rect -1518 -1150 -1506 -1116
rect -518 -1150 -506 -1116
rect -1518 -1156 -1460 -1150
rect -518 -1156 -460 -1150
rect -1518 -1328 -1460 -1322
rect -518 -1328 -460 -1322
rect -1518 -1362 -1506 -1328
rect -518 -1362 -506 -1328
rect -1518 -1368 -1460 -1362
rect -518 -1368 -460 -1362
rect -1518 -2134 -1460 -2128
rect -1018 -2134 -960 -2128
rect -518 -2134 -460 -2128
rect -1518 -2168 -1506 -2134
rect -1018 -2168 -1006 -2134
rect -518 -2168 -506 -2134
rect -1518 -2174 -1460 -2168
rect -1018 -2174 -960 -2168
rect -518 -2174 -460 -2168
rect -1518 -2328 -1460 -2322
rect -1018 -2328 -960 -2322
rect -1518 -2362 -1506 -2328
rect -1018 -2362 -1006 -2328
rect -1518 -2368 -1460 -2362
rect -1018 -2368 -960 -2362
rect -1518 -2834 -1460 -2828
rect -1518 -2868 -1506 -2834
rect -478 -2854 -420 -2848
rect -1518 -2874 -1460 -2868
rect -478 -2888 -466 -2854
rect -478 -2894 -420 -2888
<< nwell >>
rect -1416 -234 -733 -137
rect -1416 -336 -966 -234
rect -932 -336 -733 -234
rect -1416 -569 -733 -336
rect -1170 -660 -1110 -569
rect -1700 -1500 -1660 -980
<< pwell >>
rect -318 -2040 -268 -2034
rect -1340 -2450 -1130 -2040
rect -1750 -2460 -1130 -2450
rect -840 -2450 -650 -2040
rect -340 -2116 -268 -2040
rect -318 -2134 -268 -2116
rect -840 -2460 -220 -2450
rect -1750 -2760 -220 -2460
rect -1750 -3160 -1650 -2760
rect -1340 -2780 -220 -2760
rect -1340 -3160 -610 -2780
rect -290 -3160 -220 -2780
rect -1750 -3190 -220 -3160
<< psubdiff >>
rect -318 -2040 -268 -2034
rect -1340 -2450 -1130 -2040
rect -1750 -2460 -1130 -2450
rect -840 -2450 -650 -2040
rect -340 -2116 -268 -2040
rect -318 -2134 -268 -2116
rect -840 -2460 -220 -2450
rect -1750 -2760 -220 -2460
rect -1750 -3160 -1650 -2760
rect -1340 -2780 -220 -2760
rect -1340 -3160 -610 -2780
rect -290 -3160 -220 -2780
rect -1750 -3190 -220 -3160
<< locali >>
rect -2382 70 -1974 106
rect -2382 -26 -238 70
rect -2382 -108 -1652 -26
rect -468 -66 -238 -26
rect -468 -108 -240 -66
rect -2382 -234 -240 -108
rect -2382 -260 -966 -234
rect -932 -260 -240 -234
rect -2382 -320 -1100 -260
rect -2382 -660 -1110 -320
rect -966 -340 -932 -336
rect -810 -660 -240 -260
rect -2382 -1040 -240 -660
rect -2382 -1450 -1660 -1040
rect -1340 -1450 -650 -1040
rect -320 -1450 -240 -1040
rect -2382 -1498 -240 -1450
rect -2382 -1700 -238 -1498
rect -2382 -2070 -220 -1700
rect -2382 -2450 -1660 -2070
rect -1340 -2450 -1130 -2070
rect -2382 -2460 -1130 -2450
rect -840 -2450 -650 -2070
rect -340 -2116 -220 -2070
rect -320 -2450 -220 -2116
rect -840 -2460 -220 -2450
rect -2382 -2760 -220 -2460
rect -2382 -2808 -1650 -2760
rect -2382 -3144 -2046 -2808
rect -1938 -3144 -1650 -2808
rect -1340 -2780 -220 -2760
rect -2382 -3160 -1650 -3144
rect -1506 -3160 -1470 -3060
rect -1340 -3160 -610 -2780
rect -466 -3160 -432 -3048
rect -290 -3160 -220 -2780
rect -2382 -3330 -220 -3160
rect -2382 -3406 -1628 -3330
rect -328 -3406 -222 -3330
rect -2382 -3484 -222 -3406
rect -1988 -3486 -222 -3484
<< viali >>
rect -1652 -108 -468 -26
rect -2046 -3144 -1938 -2808
rect -1628 -3406 -328 -3330
<< metal1 >>
rect -3500 100 -3300 300
rect -1970 -26 -242 40
rect -1970 -108 -1652 -26
rect -468 -108 -242 -26
rect -1970 -120 -242 -108
rect -1970 -162 -240 -120
rect -1970 -164 -1770 -162
rect -966 -340 -932 -336
rect -3200 -600 -3000 -400
rect -3300 -1000 -3200 -800
rect -506 -2394 -472 -2328
rect -2110 -2808 -1840 -2560
rect -505 -2584 -473 -2394
rect -794 -2616 -473 -2584
rect -2110 -3144 -2046 -2808
rect -1938 -3144 -1840 -2808
rect -2110 -3188 -1840 -3144
rect -1506 -3264 -1470 -3060
rect -792 -3264 -763 -2616
rect -466 -3264 -432 -3048
rect -1962 -3330 -226 -3264
rect -1962 -3406 -1628 -3330
rect -328 -3406 -226 -3330
rect -1962 -3474 -226 -3406
use 10p  C1
timestamp 1742396754
transform 1 0 2900 0 1 -3374
box 0 0 1 1
use 3p  C2
timestamp 1742396754
transform 1 0 2899 0 1 -3374
box 0 0 1 1
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC1
timestamp 1742490926
transform 1 0 3006 0 1 -5040
box -3216 -3040 3216 3040
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC2
timestamp 1742490926
transform 1 0 3016 0 1 1440
box -3216 -3040 3216 3040
use sky130_fd_pr__nfet_01v8_AVVCUT  XM1
timestamp 1742490926
transform 1 0 -1489 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM2
timestamp 1742490926
transform 1 0 -989 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM3
timestamp 1742490926
transform 1 0 -1489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM4
timestamp 1742490926
transform 1 0 -489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM5
timestamp 1742490926
transform 1 0 -449 0 1 -2968
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM6
timestamp 1742490926
transform 1 0 -949 0 1 -459
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM7
timestamp 1742490926
transform 1 0 -489 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM8
timestamp 1742490926
transform 1 0 -1489 0 1 -2948
box -211 -252 211 252
<< labels >>
flabel metal1 -3500 100 -3300 300 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 -3200 -600 -3000 -400 0 FreeSans 256 0 0 0 plus
port 1 nsew
flabel metal1 -3400 -1000 -3200 -800 0 FreeSans 256 0 0 0 minus
port 0 nsew
flabel metal1 -1970 -162 -1770 38 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 -1962 -3464 -1762 -3264 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 -2080 -2770 -1880 -2570 0 FreeSans 256 0 0 0 Ibias
port 5 nsew
<< end >>
