magic
tech sky130A
magscale 1 2
timestamp 1742484632
<< checkpaint >>
rect 1692 -5058 17076 3542
<< error_s >>
rect 298 -2993 333 -2959
rect 299 -3012 333 -2993
rect 129 -3061 187 -3055
rect 129 -3095 141 -3061
rect 129 -3101 187 -3095
rect 129 -3255 187 -3249
rect 129 -3289 141 -3255
rect 129 -3295 187 -3289
rect 318 -3391 333 -3012
rect 352 -3046 387 -3012
rect 667 -3046 702 -3012
rect 352 -3391 386 -3046
rect 668 -3065 702 -3046
rect 498 -3114 556 -3108
rect 498 -3148 510 -3114
rect 498 -3154 556 -3148
rect 498 -3308 556 -3302
rect 498 -3342 510 -3308
rect 498 -3348 556 -3342
rect 352 -3425 367 -3391
rect 687 -3444 702 -3065
rect 721 -3099 756 -3065
rect 1036 -3099 1071 -3065
rect 721 -3444 755 -3099
rect 1037 -3118 1071 -3099
rect 867 -3167 925 -3161
rect 867 -3201 879 -3167
rect 867 -3207 925 -3201
rect 867 -3361 925 -3355
rect 867 -3395 879 -3361
rect 867 -3401 925 -3395
rect 721 -3478 736 -3444
rect 1056 -3497 1071 -3118
rect 1090 -3152 1125 -3118
rect 1405 -3152 1440 -3118
rect 1090 -3497 1124 -3152
rect 1406 -3171 1440 -3152
rect 1792 -3171 1845 -3170
rect 1236 -3220 1294 -3214
rect 1236 -3254 1248 -3220
rect 1236 -3260 1294 -3254
rect 1236 -3414 1294 -3408
rect 1236 -3448 1248 -3414
rect 1236 -3454 1294 -3448
rect 1090 -3531 1105 -3497
rect 1425 -3550 1440 -3171
rect 1459 -3205 1494 -3171
rect 1774 -3205 1845 -3171
rect 1459 -3550 1493 -3205
rect 1775 -3206 1845 -3205
rect 1792 -3240 1863 -3206
rect 2143 -3240 2178 -3206
rect 1605 -3273 1663 -3267
rect 1605 -3307 1617 -3273
rect 1605 -3313 1663 -3307
rect 1605 -3467 1663 -3461
rect 1605 -3501 1617 -3467
rect 1605 -3507 1663 -3501
rect 1459 -3584 1474 -3550
rect 1792 -3603 1862 -3240
rect 2144 -3259 2178 -3240
rect 1974 -3308 2032 -3302
rect 1974 -3342 1986 -3308
rect 1974 -3348 2032 -3342
rect 1974 -3520 2032 -3514
rect 1974 -3554 1986 -3520
rect 1974 -3560 2032 -3554
rect 1792 -3639 1845 -3603
rect 2163 -3656 2178 -3259
rect 2197 -3293 2232 -3259
rect 2512 -3293 2547 -3259
rect 2197 -3656 2231 -3293
rect 2513 -3312 2547 -3293
rect 2343 -3361 2401 -3355
rect 2343 -3395 2355 -3361
rect 2343 -3401 2401 -3395
rect 2343 -3573 2401 -3567
rect 2343 -3607 2355 -3573
rect 2343 -3613 2401 -3607
rect 2197 -3690 2212 -3656
rect 2532 -3709 2547 -3312
rect 2566 -3346 2601 -3312
rect 2566 -3709 2600 -3346
rect 2712 -3414 2770 -3408
rect 2712 -3448 2724 -3414
rect 2712 -3454 2770 -3448
rect 2712 -3626 2770 -3620
rect 2712 -3660 2724 -3626
rect 2712 -3666 2770 -3660
rect 2566 -3743 2581 -3709
<< pwell >>
rect 1590 -1650 1730 -1180
rect 1670 -1660 1720 -1650
rect 2040 -1680 2120 -1180
rect 1290 -1740 1330 -1680
<< locali >>
rect 670 270 1510 430
rect 670 190 2820 270
rect 670 70 970 190
rect 2690 70 2820 190
rect 670 30 2820 70
rect 680 -40 2820 30
rect 680 -440 760 -40
rect 1060 -420 1540 -40
rect 1820 -420 2460 -40
rect 1060 -440 2460 -420
rect 2760 -440 2820 -40
rect 680 -520 2820 -440
rect 720 -1240 2120 -1180
rect 720 -1640 810 -1240
rect 1130 -1640 1280 -1240
rect 1590 -1640 1730 -1240
rect 720 -1650 1730 -1640
rect 2040 -1650 2120 -1240
rect 720 -1740 2120 -1650
rect 720 -1810 930 -1740
rect 2020 -1810 2120 -1740
rect 720 -1860 2120 -1810
rect 720 -1870 1160 -1860
<< viali >>
rect 970 70 2690 190
rect 930 -1810 2020 -1740
<< metal1 >>
rect 670 260 1510 430
rect 0 0 200 200
rect 670 190 2800 260
rect 670 70 970 190
rect 2690 70 2800 190
rect 670 0 2800 70
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 720 -1740 2120 -1670
rect 0 -2000 200 -1800
rect 720 -1810 930 -1740
rect 2020 -1810 2120 -1740
rect 720 -1850 2120 -1810
rect 720 -1870 1160 -1850
use 10p  C1
timestamp 1742396754
transform 1 0 2900 0 1 -3374
box 0 0 1 1
use 3p  C2
timestamp 1742396754
transform 1 0 2899 0 1 -3374
box 0 0 1 1
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC1
timestamp 0
transform 1 0 12600 0 1 -758
box -3216 -3040 3216 3040
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC2
timestamp 0
transform 1 0 6168 0 1 -758
box -3216 -3040 3216 3040
use sky130_fd_pr__nfet_01v8_AVVCUT  XM1
timestamp 0
transform 1 0 158 0 1 -3175
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM2
timestamp 0
transform 1 0 527 0 1 -3228
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM3
timestamp 0
transform 1 0 2372 0 1 -3484
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM4
timestamp 0
transform 1 0 2003 0 1 -3431
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM5
timestamp 0
transform 1 0 896 0 1 -3281
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM6
timestamp 0
transform 1 0 2741 0 1 -3537
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM7
timestamp 0
transform 1 0 1265 0 1 -3334
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM8
timestamp 0
transform 1 0 1634 0 1 -3387
box -211 -252 211 252
<< labels >>
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 plus
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Ibias
port 5 nsew
flabel metal1 720 -1870 920 -1670 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 minus
port 0 nsew
flabel metal1 710 90 910 290 0 FreeSans 256 0 0 0 VDD
port 3 nsew
<< end >>
