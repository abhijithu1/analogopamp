magic
tech sky130A
magscale 1 2
timestamp 1742654704
<< error_s >>
rect -978 -336 -920 -330
rect -978 -370 -966 -336
rect -978 -376 -920 -370
rect -978 -548 -920 -542
rect -978 -582 -966 -548
rect -978 -588 -920 -582
rect -1518 -1116 -1460 -1110
rect -518 -1116 -460 -1110
rect -1518 -1150 -1506 -1116
rect -518 -1150 -506 -1116
rect -1518 -1156 -1460 -1150
rect -518 -1156 -460 -1150
rect -1518 -1328 -1460 -1322
rect -518 -1328 -460 -1322
rect -1518 -1362 -1506 -1328
rect -518 -1362 -506 -1328
rect -1518 -1368 -1460 -1362
rect -518 -1368 -460 -1362
rect -1518 -2328 -1460 -2322
rect -1018 -2328 -960 -2322
rect -1518 -2362 -1506 -2328
rect -1018 -2362 -1006 -2328
rect -1518 -2368 -1460 -2362
rect -1018 -2368 -960 -2362
<< nwell >>
rect -1416 -234 -733 -137
rect -1416 -336 -966 -234
rect -932 -336 -733 -234
rect -1416 -569 -733 -336
rect -1170 -660 -1110 -569
rect -1700 -1500 -1660 -980
<< pwell >>
rect -318 -2040 -268 -2034
rect -1340 -2450 -1130 -2040
rect -1750 -2460 -1130 -2450
rect -840 -2450 -650 -2040
rect -340 -2116 -268 -2040
rect -318 -2134 -268 -2116
rect -348 -2428 -286 -2270
rect -570 -2450 -286 -2428
rect -840 -2460 -220 -2450
rect -1750 -2466 -220 -2460
rect -1750 -2562 -516 -2466
rect -1750 -2630 -750 -2562
rect -1750 -2640 -516 -2630
rect -390 -2640 -220 -2466
rect -1750 -2760 -220 -2640
rect -1750 -3028 -1650 -2760
rect -1340 -2860 -220 -2760
rect -1340 -2920 -222 -2860
rect -1564 -2980 -1540 -2920
rect -1362 -2938 -222 -2920
rect -1362 -2980 -220 -2938
rect -1840 -3058 -1472 -3028
rect -1750 -3160 -1650 -3058
rect -1564 -3062 -1472 -3058
rect -1340 -3160 -220 -2980
rect -1750 -3164 -1506 -3160
rect -1470 -3162 -220 -3160
rect -1448 -3164 -220 -3162
rect -1750 -3190 -220 -3164
rect -1224 -3260 -220 -3190
rect -768 -3280 -220 -3260
rect -768 -3539 -221 -3280
<< psubdiff >>
rect -318 -2040 -268 -2034
rect -1340 -2450 -1130 -2040
rect -1750 -2460 -1130 -2450
rect -840 -2450 -650 -2040
rect -340 -2116 -268 -2040
rect -318 -2134 -268 -2116
rect -348 -2430 -286 -2270
rect -390 -2450 -286 -2430
rect -840 -2460 -516 -2450
rect -1750 -2562 -516 -2460
rect -1750 -2630 -750 -2562
rect -1750 -2640 -516 -2630
rect -390 -2640 -220 -2450
rect -1750 -2760 -220 -2640
rect -1750 -3160 -1650 -2760
rect -1340 -2780 -220 -2760
rect -1340 -2920 -610 -2780
rect -290 -2860 -220 -2780
rect -1362 -2980 -610 -2920
rect -300 -2960 -220 -2860
rect -1340 -3160 -610 -2980
rect -290 -3160 -220 -2960
rect -1750 -3164 -1506 -3160
rect -1470 -3162 -466 -3160
rect -1448 -3164 -466 -3162
rect -1750 -3184 -466 -3164
rect -432 -3184 -220 -3160
rect -1750 -3190 -220 -3184
rect -1224 -3260 -752 -3190
<< locali >>
rect -1976 106 -242 108
rect -2382 70 -242 106
rect -2382 -26 -238 70
rect -2382 -108 -1652 -26
rect -468 -66 -238 -26
rect -468 -108 -240 -66
rect -2382 -234 -240 -108
rect -2382 -260 -966 -234
rect -932 -260 -240 -234
rect -2382 -320 -1100 -260
rect -2382 -660 -1110 -320
rect -966 -340 -932 -336
rect -810 -660 -240 -260
rect -2382 -1040 -240 -660
rect -2382 -1450 -1660 -1040
rect -1340 -1450 -650 -1040
rect -320 -1450 -240 -1040
rect -2382 -1498 -240 -1450
rect -2382 -1580 -238 -1498
rect -2382 -1656 -2170 -1580
rect -1740 -1656 -238 -1580
rect -2382 -1700 -238 -1656
rect -2382 -2012 -220 -1700
rect -2382 -2422 -2248 -2012
rect -2126 -2070 -220 -2012
rect -2126 -2422 -1660 -2070
rect -2382 -2450 -1660 -2422
rect -1340 -2450 -1130 -2070
rect -2382 -2460 -1130 -2450
rect -840 -2450 -650 -2070
rect -340 -2116 -220 -2070
rect -320 -2270 -220 -2116
rect -348 -2430 -220 -2270
rect -516 -2450 -220 -2430
rect -840 -2460 -220 -2450
rect -2382 -2760 -220 -2460
rect -2382 -2808 -1650 -2760
rect -2382 -3144 -2046 -2808
rect -1938 -2920 -1650 -2808
rect -1340 -2780 -220 -2760
rect -1340 -2920 -610 -2780
rect -1938 -2980 -1540 -2920
rect -1362 -2980 -610 -2920
rect -1938 -3028 -1650 -2980
rect -1938 -3060 -1472 -3028
rect -1938 -3062 -1470 -3060
rect -1938 -3144 -1650 -3062
rect -1506 -3068 -1470 -3062
rect -2382 -3160 -1650 -3144
rect -1506 -3156 -1470 -3130
rect -1506 -3158 -1444 -3156
rect -1506 -3160 -1438 -3158
rect -1340 -3160 -610 -2980
rect -466 -3082 -432 -3048
rect -528 -3160 -370 -3150
rect -300 -3160 -220 -2780
rect -2382 -3162 -220 -3160
rect -2382 -3164 -1474 -3162
rect -1448 -3164 -220 -3162
rect -2382 -3330 -220 -3164
rect -2382 -3406 -1628 -3330
rect -328 -3406 -222 -3330
rect -2382 -3484 -222 -3406
rect -1988 -3486 -222 -3484
<< viali >>
rect -1652 -108 -468 -26
rect -2170 -1656 -1740 -1580
rect -2248 -2422 -2126 -2012
rect -2046 -3144 -1938 -2808
rect -1628 -3406 -328 -3330
<< metal1 >>
rect -3500 100 -3300 300
rect -1970 -26 -242 40
rect -1970 -108 -1652 -26
rect -468 -108 -242 -26
rect -1970 -120 -242 -108
rect -1970 -162 -240 -120
rect -1970 -164 -1770 -162
rect -966 -340 -932 -336
rect -2378 -1580 -1712 -1538
rect -2378 -1656 -2170 -1580
rect -1740 -1656 -1712 -1580
rect -2378 -1738 -1712 -1656
rect -2178 -1740 -1712 -1738
rect -2302 -2012 -2048 -1778
rect -2302 -2422 -2248 -2012
rect -2126 -2422 -2048 -2012
rect -428 -2278 -286 -2218
rect -1506 -2362 -1472 -2328
rect -506 -2333 -472 -2328
rect -703 -2362 -472 -2333
rect -2302 -2474 -2048 -2422
rect -703 -2363 -503 -2362
rect -1570 -2466 -910 -2430
rect -2110 -2642 -1840 -2560
rect -703 -2642 -673 -2363
rect -348 -2428 -286 -2278
rect -570 -2466 -286 -2428
rect -2110 -2672 -673 -2642
rect -390 -2468 -286 -2466
rect -390 -2582 -314 -2468
rect -390 -2584 -262 -2582
rect -390 -2652 -220 -2584
rect -2110 -2808 -1840 -2672
rect -2110 -3144 -2046 -2808
rect -1938 -2920 -1840 -2808
rect -1462 -2920 -1360 -2918
rect -1938 -2980 -1540 -2920
rect -1462 -2980 -1224 -2920
rect -1938 -3028 -1840 -2980
rect -1938 -3060 -1472 -3028
rect -1938 -3062 -1470 -3060
rect -1938 -3144 -1840 -3062
rect -2110 -3188 -1840 -3144
rect -1568 -3142 -1410 -3130
rect -1274 -3142 -1224 -2980
rect -703 -3050 -673 -2672
rect -300 -2938 -220 -2652
rect -406 -2996 -220 -2938
rect -630 -3050 -432 -3048
rect -703 -3079 -432 -3050
rect -700 -3080 -432 -3079
rect -466 -3082 -432 -3080
rect -1568 -3202 -1224 -3142
rect -792 -3264 -763 -3260
rect -528 -3264 -370 -3150
rect -300 -3264 -220 -2996
rect -1962 -3280 -220 -3264
rect -1962 -3330 -226 -3280
rect -1962 -3406 -1628 -3330
rect -328 -3406 -226 -3330
rect -1962 -3474 -226 -3406
use 10p  C1
timestamp 1742396754
transform 1 0 2900 0 1 -3374
box 0 0 1 1
use 3p  C2
timestamp 1742396754
transform 1 0 2899 0 1 -3374
box 0 0 1 1
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC1
timestamp 1742490926
transform 1 0 3006 0 1 -5040
box -3216 -3040 3216 3040
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC2
timestamp 1742490926
transform 1 0 3016 0 1 1440
box -3216 -3040 3216 3040
use sky130_fd_pr__nfet_01v8_AVVCUT  XM1
timestamp 1742648969
transform 1 0 -1489 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM2
timestamp 1742648969
transform 1 0 -989 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM3
timestamp 1742490926
transform 1 0 -1489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM4
timestamp 1742490926
transform 1 0 -489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM5
timestamp 1742648969
transform 1 0 -449 0 1 -2968
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM6
timestamp 1742490926
transform 1 0 -949 0 1 -459
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM7
timestamp 1742648969
transform 1 0 -489 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM8
timestamp 1742648969
transform 1 0 -1489 0 1 -2948
box -211 -252 211 252
<< labels >>
flabel metal1 -3500 100 -3300 300 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 -1970 -162 -1770 38 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 -1962 -3464 -1762 -3264 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 -2080 -2770 -1880 -2570 0 FreeSans 256 0 0 0 Ibias
port 5 nsew
flabel metal1 -2278 -1988 -2078 -1788 0 FreeSans 256 0 0 0 plus
port 1 nsew
flabel metal1 -2378 -1738 -2178 -1538 0 FreeSans 256 0 0 0 minus
port 0 nsew
<< end >>
