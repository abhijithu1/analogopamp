magic
tech sky130A
magscale 1 2
timestamp 1742490926
<< error_s >>
rect -978 -336 -920 -330
rect -978 -370 -966 -336
rect -978 -376 -920 -370
rect -978 -548 -920 -542
rect -978 -582 -966 -548
rect -978 -588 -920 -582
rect -1518 -1116 -1460 -1110
rect -518 -1116 -460 -1110
rect -1518 -1150 -1506 -1116
rect -518 -1150 -506 -1116
rect -1518 -1156 -1460 -1150
rect -518 -1156 -460 -1150
rect -1518 -1328 -1460 -1322
rect -518 -1328 -460 -1322
rect -1518 -1362 -1506 -1328
rect -518 -1362 -506 -1328
rect -1518 -1368 -1460 -1362
rect -518 -1368 -460 -1362
rect -1518 -2134 -1460 -2128
rect -1018 -2134 -960 -2128
rect -518 -2134 -460 -2128
rect -1518 -2168 -1506 -2134
rect -1018 -2168 -1006 -2134
rect -518 -2168 -506 -2134
rect -1518 -2174 -1460 -2168
rect -1018 -2174 -960 -2168
rect -518 -2174 -460 -2168
rect -1518 -2328 -1460 -2322
rect -1018 -2328 -960 -2322
rect -518 -2328 -460 -2322
rect -1518 -2362 -1506 -2328
rect -1018 -2362 -1006 -2328
rect -518 -2362 -506 -2328
rect -1518 -2368 -1460 -2362
rect -1018 -2368 -960 -2362
rect -518 -2368 -460 -2362
rect -1518 -2834 -1460 -2828
rect -1518 -2868 -1506 -2834
rect -478 -2854 -420 -2848
rect -1518 -2874 -1460 -2868
rect -478 -2888 -466 -2854
rect -478 -2894 -420 -2888
rect -1518 -3028 -1460 -3022
rect -1518 -3062 -1506 -3028
rect -478 -3048 -420 -3042
rect -1518 -3068 -1460 -3062
rect -478 -3082 -466 -3048
rect -478 -3088 -420 -3082
<< nwell >>
rect -1170 -260 -740 -180
rect -1170 -320 -1100 -260
rect -1170 -660 -1110 -320
rect -1700 -1500 -1660 -980
<< pwell >>
rect -1340 -2450 -1130 -2040
rect -1750 -2460 -1130 -2450
rect -840 -2450 -650 -2040
rect -840 -2460 -220 -2450
rect -1750 -2760 -220 -2460
rect -1750 -3160 -1650 -2760
rect -1340 -2780 -220 -2760
rect -1340 -3160 -610 -2780
rect -290 -3160 -220 -2780
rect -1750 -3190 -220 -3160
<< psubdiff >>
rect -1340 -2450 -1130 -2040
rect -1750 -2460 -1130 -2450
rect -840 -2450 -650 -2040
rect -840 -2460 -220 -2450
rect -1750 -2760 -220 -2460
rect -1750 -3160 -1650 -2760
rect -1340 -2780 -220 -2760
rect -1340 -3160 -610 -2780
rect -290 -3160 -220 -2780
rect -1750 -3190 -220 -3160
<< locali >>
rect -1710 -80 -240 -50
rect -1710 -160 -1610 -80
rect -410 -160 -240 -80
rect -1710 -260 -240 -160
rect -1710 -320 -1100 -260
rect -1710 -660 -1110 -320
rect -810 -660 -240 -260
rect -1710 -1000 -240 -660
rect -1700 -1040 -240 -1000
rect -1700 -1450 -1660 -1040
rect -1340 -1450 -650 -1040
rect -320 -1450 -240 -1040
rect -1700 -1510 -240 -1450
rect -1750 -2070 -220 -1700
rect -1750 -2450 -1660 -2070
rect -1340 -2450 -1130 -2070
rect -1750 -2460 -1130 -2450
rect -840 -2450 -650 -2070
rect -320 -2450 -220 -2070
rect -840 -2460 -220 -2450
rect -1750 -2760 -220 -2460
rect -1750 -3160 -1650 -2760
rect -1340 -2780 -220 -2760
rect -1340 -3160 -610 -2780
rect -290 -3160 -220 -2780
rect -1750 -3230 -220 -3160
rect -1750 -3300 -1640 -3230
rect -320 -3300 -220 -3230
rect -1750 -3330 -220 -3300
<< viali >>
rect -1610 -160 -410 -80
rect -1640 -3300 -320 -3230
<< metal1 >>
rect -3500 100 -3300 300
rect -3500 -200 -3300 0
rect -1700 -80 -280 -70
rect -1700 -160 -1610 -80
rect -410 -160 -280 -80
rect -1700 -170 -280 -160
rect -3500 -500 -3300 -300
rect -3200 -600 -3000 -400
rect -3400 -1000 -3200 -800
rect -3500 -1400 -3300 -1196
rect -1730 -3230 -250 -3200
rect -1730 -3300 -1640 -3230
rect -320 -3300 -250 -3230
rect -1730 -3330 -250 -3300
use 10p  C1
timestamp 1742396754
transform 1 0 2900 0 1 -3374
box 0 0 1 1
use 3p  C2
timestamp 1742396754
transform 1 0 2899 0 1 -3374
box 0 0 1 1
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC1
timestamp 1742490926
transform 1 0 3006 0 1 -5040
box -3216 -3040 3216 3040
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC2
timestamp 1742490926
transform 1 0 3016 0 1 1440
box -3216 -3040 3216 3040
use sky130_fd_pr__nfet_01v8_AVVCUT  XM1
timestamp 1742490926
transform 1 0 -1489 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM2
timestamp 1742490926
transform 1 0 -989 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM3
timestamp 1742490926
transform 1 0 -1489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM4
timestamp 1742490926
transform 1 0 -489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM5
timestamp 1742490926
transform 1 0 -449 0 1 -2968
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM6
timestamp 1742490926
transform 1 0 -949 0 1 -459
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM7
timestamp 1742490926
transform 1 0 -489 0 1 -2248
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM8
timestamp 1742490926
transform 1 0 -1489 0 1 -2948
box -211 -252 211 252
<< labels >>
flabel metal1 -3500 100 -3300 300 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 -3500 -200 -3300 0 0 FreeSans 256 0 0 0 Ibias
port 5 nsew
flabel metal1 -3500 -500 -3300 -300 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 -3200 -600 -3000 -400 0 FreeSans 256 0 0 0 plus
port 1 nsew
flabel metal1 -3400 -1000 -3200 -800 0 FreeSans 256 0 0 0 minus
port 0 nsew
flabel metal1 -3500 -1398 -3300 -1198 0 FreeSans 256 0 0 0 VDD
port 3 nsew
<< end >>
