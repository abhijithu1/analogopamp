magic
tech sky130A
timestamp 1742396754
<< end >>
