magic
tech sky130A
magscale 1 2
timestamp 1742985680
<< nwell >>
rect -1170 -260 -740 -180
rect -1170 -320 -1100 -260
rect -1170 -660 -1110 -320
rect -1700 -1500 -1660 -980
rect -1506 -1120 -1282 -1116
rect -1278 -1120 -1276 -1042
rect -1506 -1122 -1276 -1120
rect -1506 -1150 -1292 -1122
rect -1310 -1210 -1292 -1150
rect -1282 -1210 -1276 -1122
rect -622 -1150 -548 -1102
rect -1310 -1216 -1284 -1210
<< pwell >>
rect -1272 -1268 -1166 -1210
rect -2532 -1540 -2462 -1538
rect -1230 -1540 -1166 -1268
rect -2532 -1610 -1166 -1540
rect -2790 -2288 -2692 -2054
rect -2532 -2180 -2462 -1610
rect -712 -1878 -650 -1876
rect -1962 -1880 -648 -1878
rect -1964 -1934 -648 -1880
rect -1964 -2180 -1896 -1934
rect -2532 -2238 -2278 -2180
rect -2532 -2242 -2462 -2238
rect -2224 -2240 -1894 -2180
rect -1582 -2288 -1412 -1980
rect -712 -2180 -650 -1934
rect -914 -2240 -650 -2180
rect -712 -2242 -650 -2240
rect 150 -2286 186 -2174
rect 388 -2246 688 -2186
rect -2790 -2290 -2466 -2288
rect -1582 -2290 -1168 -2288
rect -2790 -2324 -2234 -2290
rect -1582 -2322 -924 -2290
rect -2790 -2412 -2692 -2324
rect -2330 -2498 -2174 -2372
rect -1582 -2456 -1412 -2322
rect -1218 -2324 -924 -2322
rect 250 -2330 290 -2296
rect -1020 -2468 -862 -2374
rect -974 -2498 -908 -2468
rect -2330 -2562 -908 -2498
rect -2330 -2566 -954 -2562
rect -2330 -2568 -2174 -2566
rect -1910 -2568 -1574 -2566
rect -402 -3378 -82 -3318
<< locali >>
rect -2926 8096 3672 8118
rect -2926 5736 13864 8096
rect -2926 1876 3672 5736
rect -2926 1702 3704 1876
rect -2896 1422 3704 1702
rect -2896 1174 -1422 1422
rect 1348 1174 3704 1422
rect -2896 398 3704 1174
rect -2900 -178 3704 398
rect -2898 -252 3704 -178
rect 10090 -210 13830 5736
rect 10062 -252 13830 -210
rect -2898 -258 13830 -252
rect -2898 -260 13818 -258
rect -2898 -320 -1100 -260
rect -1028 -274 -866 -260
rect -2898 -428 -1110 -320
rect -810 -336 13818 -260
rect -966 -370 13818 -336
rect -2898 -488 -976 -428
rect -2898 -660 -1110 -488
rect -810 -660 13818 -370
rect -2898 -1040 13818 -660
rect -2898 -1450 -1660 -1040
rect -1566 -1078 -1410 -1040
rect -1340 -1114 -650 -1040
rect -1356 -1150 -650 -1114
rect -1340 -1450 -650 -1150
rect -320 -1208 13818 -1040
rect -462 -1270 13818 -1208
rect -320 -1450 13818 -1270
rect -2898 -1454 13818 -1450
rect -2912 -1534 13818 -1454
rect -2912 -2014 3646 -1534
rect -2910 -2180 -2408 -2014
rect -2090 -2180 -1098 -2014
rect -784 -2180 214 -2014
rect -2910 -2192 -2278 -2180
rect -2910 -2400 -2776 -2192
rect -2726 -2238 -2278 -2192
rect -2224 -2200 -968 -2180
rect -2726 -2290 -2408 -2238
rect -2224 -2240 -1556 -2200
rect -2726 -2324 -2234 -2290
rect -2726 -2400 -2408 -2324
rect -2910 -2416 -2408 -2400
rect -2330 -2416 -2174 -2372
rect -2090 -2416 -1556 -2240
rect -2914 -2430 -1556 -2416
rect -1452 -2238 -968 -2200
rect -914 -2186 214 -2180
rect 526 -2186 3646 -2014
rect -1452 -2290 -1098 -2238
rect -914 -2240 334 -2186
rect -784 -2246 334 -2240
rect 388 -2246 3646 -2186
rect -1452 -2324 -924 -2290
rect -784 -2296 214 -2246
rect -1452 -2416 -1098 -2324
rect -784 -2330 276 -2296
rect -1020 -2416 -862 -2374
rect -784 -2416 214 -2330
rect 282 -2416 448 -2398
rect 526 -2416 3646 -2246
rect -1452 -2430 3646 -2416
rect -2914 -2486 3646 -2430
rect -2932 -2702 3646 -2486
rect -2934 -3150 3646 -2702
rect -2934 -3310 -1740 -3150
rect -2934 -3336 -1610 -3310
rect -2934 -3548 -2218 -3336
rect -2158 -3374 -1610 -3336
rect -2158 -3422 -1740 -3374
rect -2158 -3456 -1566 -3422
rect -1424 -3428 -582 -3150
rect -270 -3318 3646 -3150
rect -402 -3378 3646 -3318
rect -2158 -3542 -1740 -3456
rect -1424 -3462 -410 -3428
rect -1664 -3542 -1506 -3506
rect -1424 -3542 -582 -3462
rect -2158 -3548 -582 -3542
rect -2934 -3552 -582 -3548
rect -512 -3552 -344 -3508
rect -270 -3552 3646 -3378
rect -2934 -3942 3646 -3552
rect -2938 -4752 3646 -3942
rect -2938 -4968 -1532 -4752
rect 1412 -4968 3646 -4752
rect -2938 -5164 3646 -4968
rect -2934 -7576 3646 -5164
rect 10062 -7482 13818 -1534
rect 10060 -7562 13818 -7482
rect 10060 -7574 13808 -7562
rect 9852 -7576 13808 -7574
rect -2950 -8776 13808 -7576
rect -2950 -11328 13806 -8776
<< viali >>
rect -1422 1174 1348 1422
rect -2776 -2400 -2726 -2192
rect -1556 -2430 -1452 -2200
rect -2218 -3548 -2158 -3336
rect -1532 -4968 1412 -4752
<< metal1 >>
rect -2812 1422 1476 1466
rect -2812 1174 -1422 1422
rect 1348 1174 1476 1422
rect -2812 904 1476 1174
rect -1796 -844 -1730 904
rect -1290 -18 -1222 -16
rect -980 -18 -914 904
rect -1290 -86 -866 -18
rect -1290 -428 -1222 -86
rect -1028 -274 -866 -86
rect -576 -336 -408 904
rect 1908 -310 1918 -256
rect -226 -314 1918 -310
rect -328 -336 -308 -314
rect -966 -370 -730 -336
rect -576 -372 -308 -336
rect -242 -372 1918 -314
rect -1292 -488 -976 -428
rect -1522 -844 -1452 -842
rect -1796 -896 -1410 -844
rect -1796 -1210 -1730 -896
rect -1566 -1078 -1410 -896
rect -806 -862 -740 -860
rect -576 -862 -408 -372
rect -200 -750 -144 -372
rect 1908 -416 1918 -372
rect 2368 -416 2378 -256
rect -200 -792 -142 -750
rect -806 -934 -408 -862
rect -1036 -1114 -1026 -1098
rect -1356 -1116 -1026 -1114
rect -1506 -1150 -1026 -1116
rect -974 -1150 -964 -1098
rect -1310 -1210 -1282 -1150
rect -806 -1208 -740 -934
rect -570 -1070 -408 -934
rect -484 -1072 -408 -1070
rect -632 -1150 -622 -1098
rect -570 -1102 -560 -1098
rect -570 -1116 -548 -1102
rect -570 -1150 -472 -1116
rect -198 -1208 -142 -792
rect -1796 -1270 -1516 -1210
rect -1462 -1268 -1166 -1210
rect -1796 -1272 -1730 -1270
rect -2532 -1540 -2462 -1538
rect -1230 -1540 -1166 -1268
rect -806 -1268 -514 -1208
rect -208 -1264 -198 -1208
rect -144 -1264 -134 -1208
rect -806 -1272 -740 -1268
rect -2532 -1610 -1166 -1540
rect -2836 -2096 -2636 -1896
rect -2790 -2192 -2692 -2096
rect -2790 -2400 -2776 -2192
rect -2726 -2288 -2692 -2192
rect -2532 -2180 -2462 -1610
rect 1292 -1780 1492 -1710
rect 1076 -1792 1492 -1780
rect 1076 -1844 1118 -1792
rect 1170 -1844 1492 -1792
rect 1076 -1864 1492 -1844
rect -712 -1878 -650 -1876
rect -1962 -1880 -648 -1878
rect -1964 -1934 -648 -1880
rect 1292 -1910 1492 -1864
rect -1964 -2180 -1896 -1934
rect -1440 -2000 -1412 -1980
rect -2532 -2238 -2278 -2180
rect -2532 -2242 -2462 -2238
rect -2224 -2240 -1894 -2180
rect -1592 -2200 -1392 -2000
rect -712 -2180 -650 -1934
rect -914 -2182 -650 -2180
rect -2726 -2290 -2466 -2288
rect -2726 -2324 -2234 -2290
rect -2726 -2400 -2692 -2324
rect -2790 -2412 -2692 -2400
rect -2330 -2498 -2174 -2372
rect -1582 -2430 -1556 -2200
rect -1452 -2288 -1412 -2200
rect -914 -2240 -734 -2182
rect -664 -2240 -650 -2182
rect -712 -2242 -650 -2240
rect 388 -2246 688 -2186
rect -1452 -2290 -1168 -2288
rect -1452 -2322 -924 -2290
rect -1452 -2430 -1412 -2322
rect -1218 -2324 -924 -2322
rect 260 -2330 378 -2296
rect -1582 -2456 -1412 -2430
rect -1020 -2496 -862 -2374
rect 282 -2462 448 -2398
rect 624 -2462 688 -2246
rect 282 -2496 688 -2462
rect -1020 -2498 688 -2496
rect -2330 -2514 688 -2498
rect -2330 -2562 448 -2514
rect -2330 -2564 398 -2562
rect -2330 -2566 -954 -2564
rect -2330 -2568 -2174 -2566
rect -1910 -2568 -1574 -2566
rect -220 -2912 -80 -2910
rect -860 -2914 -80 -2912
rect -1890 -2968 -80 -2914
rect -2284 -3192 -2084 -2992
rect -1890 -3028 -1844 -2968
rect -860 -2972 -80 -2968
rect -1892 -3100 -1844 -3028
rect -2236 -3310 -2132 -3192
rect -1892 -3310 -1846 -3100
rect -2236 -3336 -1610 -3310
rect -2236 -3548 -2218 -3336
rect -2158 -3372 -1610 -3336
rect -1558 -3372 -1296 -3312
rect -2158 -3548 -2132 -3372
rect -1892 -3374 -1610 -3372
rect -1892 -3422 -1846 -3374
rect -1892 -3456 -1566 -3422
rect -1892 -3460 -1846 -3456
rect -2236 -3566 -2132 -3548
rect -1664 -3578 -1506 -3506
rect -1356 -3578 -1296 -3372
rect -858 -3428 -786 -2972
rect -112 -2974 -80 -2972
rect 10 -2974 20 -2910
rect 330 -3130 398 -2564
rect -402 -3378 -82 -3318
rect -858 -3462 -410 -3428
rect -858 -3464 -786 -3462
rect -1664 -3626 -1296 -3578
rect -512 -3578 -344 -3508
rect -142 -3578 -82 -3378
rect -1664 -4620 -1506 -3626
rect -512 -3630 -82 -3578
rect -512 -4620 -344 -3630
rect 326 -4620 398 -3130
rect -2890 -4664 1596 -4620
rect -2892 -4752 1596 -4664
rect -2892 -4968 -1532 -4752
rect 1412 -4968 1596 -4752
rect -2892 -4990 1596 -4968
rect -2890 -5100 1596 -4990
<< via1 >>
rect -308 -372 -242 -314
rect 1918 -416 2368 -256
rect -1026 -1150 -974 -1098
rect -622 -1150 -570 -1098
rect -198 -1264 -144 -1208
rect 1118 -1844 1170 -1792
rect -734 -2240 -664 -2182
rect -80 -2974 10 -2910
<< metal2 >>
rect 1918 -256 2368 -246
rect -308 -314 -242 -304
rect -328 -336 -308 -314
rect -762 -370 -308 -336
rect -454 -372 -308 -370
rect -308 -382 -242 -372
rect 2368 -416 2370 -256
rect 1918 -426 2368 -416
rect -922 -488 124 -428
rect -1026 -1098 -974 -1088
rect -622 -1098 -570 -1088
rect -974 -1150 -622 -1102
rect -570 -1150 -564 -1102
rect -1026 -1160 -974 -1150
rect -622 -1160 -570 -1150
rect -198 -1208 -144 -1198
rect -462 -1264 -198 -1208
rect -144 -1264 -118 -1208
rect -462 -1270 -118 -1264
rect -198 -1274 -118 -1270
rect -178 -1728 -118 -1274
rect -1272 -1780 -118 -1728
rect 60 -1780 124 -488
rect -1272 -1854 -1206 -1780
rect 56 -1792 1202 -1780
rect 56 -1844 1118 -1792
rect 1170 -1844 1202 -1792
rect -1272 -2180 -1208 -1854
rect 56 -1862 1202 -1844
rect 60 -2008 124 -1862
rect -1272 -2238 -968 -2180
rect -734 -2182 -664 -2172
rect -1272 -2240 -1208 -2238
rect -734 -2828 -664 -2240
rect 62 -2186 124 -2008
rect 62 -2246 334 -2186
rect -80 -2296 8 -2294
rect -80 -2330 276 -2296
rect -80 -2558 8 -2330
rect -734 -3316 -666 -2828
rect -80 -2910 10 -2558
rect -80 -2984 10 -2974
rect -736 -3378 -456 -3316
<< via2 >>
rect 1918 -416 2368 -256
<< metal3 >>
rect 1908 -256 2378 -251
rect 1908 -416 1918 -256
rect 2368 -416 2378 -256
rect 1908 -421 2378 -416
<< via3 >>
rect 1926 -414 2368 -256
<< metal4 >>
rect 1930 6588 2346 6592
rect 5960 6588 12054 6594
rect 1508 6582 12054 6588
rect 1508 6126 12066 6582
rect 1508 6120 6118 6126
rect 1930 2602 2346 6120
rect 11452 4272 12066 6126
rect 10020 3646 12066 4272
rect 11452 3640 12066 3646
rect 1930 122 2358 2602
rect 1928 -255 2368 122
rect 1925 -256 2369 -255
rect 1925 -414 1926 -256
rect 2368 -414 2369 -256
rect 1925 -415 2369 -414
use 10p  C1
timestamp 1742396754
transform 1 0 2900 0 1 -3374
box 0 0 1 1
use 3p  C2
timestamp 1742396754
transform 1 0 2899 0 1 -3374
box 0 0 1 1
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC1
timestamp 1742490926
transform 1 0 6842 0 1 -4542
box -3216 -3040 3216 3040
use sky130_fd_pr__cap_mim_m3_1_8WUMYD  XC2
timestamp 1742490926
transform 1 0 6888 0 1 2750
box -3216 -3040 3216 3040
use sky130_fd_pr__nfet_01v8_AVVCUT  XM1
timestamp 1742907183
transform 1 0 -2251 0 1 -2210
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM2
timestamp 1742907183
transform 1 0 -941 0 1 -2210
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM3
timestamp 1742907183
transform 1 0 -1489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM4
timestamp 1742907183
transform 1 0 -489 0 1 -1239
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM5
timestamp 1742907183
transform 1 0 -429 0 1 -3348
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_Q3HK3C  XM6
timestamp 1742907183
transform 1 0 -949 0 1 -459
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_AVVCUT  XM7
timestamp 1742907183
transform 1 0 361 0 1 -2216
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_AVVCUT  XM8
timestamp 1742907183
transform 1 0 -1585 0 1 -3342
box -211 -252 211 252
<< labels >>
flabel metal1 -2590 1104 -2390 1304 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 -2728 -4960 -2528 -4760 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 -2836 -2096 -2636 -1896 0 FreeSans 256 0 0 0 minus
port 0 nsew
flabel metal1 -1592 -2200 -1392 -2000 0 FreeSans 256 0 0 0 plus
port 1 nsew
flabel metal1 -2284 -3192 -2084 -2992 0 FreeSans 256 0 0 0 Ibias
port 5 nsew
flabel metal1 1292 -1910 1492 -1710 0 FreeSans 256 0 0 0 Vout
port 2 nsew
<< end >>
